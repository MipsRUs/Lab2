module processor_tb;
	
  timeunit 1ns;

  logic ref_clk;
  logic reset;
  
processor L1(
          .ref_clk(ref_clk)
         ,.reset(reset)
         );

always begin
	#5 ref_clk = 1;
	#5 ref_clk = 0;
end

initial begin

	reset = 1;
	#20;
	reset = 0;
	#2000;


end
endmodule
    
